//////////////////////////////////////////////////////////////////////////////////
// File Name: 		AHB_mux.sv
// Project Name:	AHB_Gen
// Email:         quanghungbk1999@gmail.com
// Version    Date      Author      Description
// v0.0       2/10/2020 Quang Hung  First Creation
//////////////////////////////////////////////////////////////////////////////////

import AHB_package::*;
module AHB_bus
#(
  parameter AHB
)
(

);


endmodule: AHB_bus
