/*********************************************************************************
 * File Name: 		AHB_coverage.sv
 * Project Name:	AHB_Gen
 * Email:         quanghungbk1999@gmail.com
 * Version    Date       Author      Description
 * v0.0       02/10/2020 Quang Hung  First Creation
 *            12/01/2021 Quang Hung  Add support for decode error
 *            12/01/2021 Quang Hung  Config maximum cells per masters
 *            16/01/2021 Quang Hung  Add coverage support
 *********************************************************************************/

class Mas_coverage

endclass: Mas_coverage

class Slv_coverage

endclass: Slv_coverage
