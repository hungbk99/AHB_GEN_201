//////////////////////////////////////////////////////////////////////////////////
// File Name: 		arbiter_package.sv
// Project Name:	AHB_Gen
// Email:         quanghungbk1999@gmail.com
// Version    Date      Author      Description
// v0.0       9/10/2020 Quang Hung  First Creation
//////////////////////////////////////////////////////////////////////////////////

package arbiter_package;
  parameter SLAVE_0_PRIOR_NUM = 4;
  parameter SLAVE_0_PRIOR_BIT =2;
  parameter SLAVE_0_MASTER_NUM = 10;  

endpackage
